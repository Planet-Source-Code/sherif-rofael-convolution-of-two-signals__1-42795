If LengthA > LengthB Then
        Ref = LengthA
        InvRef = LengthB
    Else
        Ref = LengthB
        InvRef = LengthA
        MatrixB = Middle
        MatrixB = MatrixA
        MatrixA = Middle
    End If