Convolution of Two input signals by sherif rofael ,  First Time in planet source code , advanced code ,

